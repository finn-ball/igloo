`ifndef TOP_SIM_VH

 `define TOP_SIM_VH

 `timescale 1ns/1ps
 `define SIM 1

`endif
