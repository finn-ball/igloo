`ifndef UART_VH

 `define UART_VH

 `define UART_CLK_PERIOD 625
 `define UART_DATA_WIDTH 8

`endif
