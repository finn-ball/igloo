`include "uart.vh"

module uart_ctrl(
		 input 				   clk_i,
		 output [`UART_DATA_WIDTH - 1 : 0] tx,
		 output 			   tx_v
		 );


   
endmodule // uart_ctrl
