`include "uart.vh"

module uart_ctrl(
		 input clk_i
		 );


endmodule // uart_ctrl
