`ifndef UART_VH
 `define UART_VH

`define UART_ADDR_WIDTH 4

`endif
