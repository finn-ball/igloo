`ifndef UART_VH

 `define UART_VH

 `define UART_RX_SAMPLE_RATE 16 // NOTE, make it a power of 2
 `define UART_CLK_RX_PERIOD 625 
 `define UART_CLK_TX_PERIOD 625

 `define UART_DATA_WIDTH 8

`endif
